/********
seqDetect_tb.sv

Written by Jimmy Bates (A01035957)

ELEX 7660-Digital System Design
Assignment 2

Date created: February 12, 2022

Test bench for sequence detector

code for modelsim:
vsim work.seqDetect_tb; add wave sim:*; run -all

*********/

//Instantiate model

//Reset

//Round 1
//Store some set of bits in a 6 bit word
//Setup correct input
//Run clock 9 times

//Reset

//Round 2
//Store some set of bits in a 6 bit word
//Set up correct input
//Run clock 9 times

//stop